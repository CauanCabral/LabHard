entity barrel_shifter is
	port(
		din1, din2, din3, din4: in bit;
		desloc1, desloc2: in bit;
		dout1, dout2, dout3, dout4: out bit;
	);
end entity;


